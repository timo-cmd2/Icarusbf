`default_nettype none

module ibf
endmodule

module ibf
